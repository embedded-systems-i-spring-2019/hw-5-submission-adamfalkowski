library IEEE;
use IEEE.std_logic_1164.all;

entity crk2 is
  port (
        A_1, A_2, B_1, B_2, D_1 : in std_logic;
	      E_out : out std_logic
       );
 end crk2;
 
 architecture if_arc of crk2 
 
 
